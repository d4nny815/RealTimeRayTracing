import Primitives::*;

module TransformModule (
    input Face_t

    );


endmodule