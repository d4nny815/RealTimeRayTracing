

module GPU (



    );


    localparam FACES = 92;
    logic [$clog2(FACES) - 1 : 0] face_cntr;



endmodule