module ProjectionModule (
    

    );


endmodule